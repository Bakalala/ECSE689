-- FSM Controller
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity Controller is
    Port ( clk, rst : in STD_LOGIC;
           R0_en : out STD_LOGIC;
           R1_en : out STD_LOGIC;
           R10_en : out STD_LOGIC;
           R11_en : out STD_LOGIC;
           R12_en : out STD_LOGIC;
           R13_en : out STD_LOGIC;
           R14_en : out STD_LOGIC;
           R15_en : out STD_LOGIC;
           R16_en : out STD_LOGIC;
           R17_en : out STD_LOGIC;
           R18_en : out STD_LOGIC;
           R19_en : out STD_LOGIC;
           R2_en : out STD_LOGIC;
           R20_en : out STD_LOGIC;
           R21_en : out STD_LOGIC;
           R22_en : out STD_LOGIC;
           R23_en : out STD_LOGIC;
           R24_en : out STD_LOGIC;
           R25_en : out STD_LOGIC;
           R26_en : out STD_LOGIC;
           R27_en : out STD_LOGIC;
           R28_en : out STD_LOGIC;
           R29_en : out STD_LOGIC;
           R3_en : out STD_LOGIC;
           R30_en : out STD_LOGIC;
           R31_en : out STD_LOGIC;
           R32_en : out STD_LOGIC;
           R33_en : out STD_LOGIC;
           R34_en : out STD_LOGIC;
           R35_en : out STD_LOGIC;
           R36_en : out STD_LOGIC;
           R37_en : out STD_LOGIC;
           R38_en : out STD_LOGIC;
           R39_en : out STD_LOGIC;
           R4_en : out STD_LOGIC;
           R40_en : out STD_LOGIC;
           R41_en : out STD_LOGIC;
           R42_en : out STD_LOGIC;
           R43_en : out STD_LOGIC;
           R44_en : out STD_LOGIC;
           R45_en : out STD_LOGIC;
           R46_en : out STD_LOGIC;
           R47_en : out STD_LOGIC;
           R48_en : out STD_LOGIC;
           R49_en : out STD_LOGIC;
           R5_en : out STD_LOGIC;
           R50_en : out STD_LOGIC;
           R51_en : out STD_LOGIC;
           R52_en : out STD_LOGIC;
           R53_en : out STD_LOGIC;
           R54_en : out STD_LOGIC;
           R55_en : out STD_LOGIC;
           R56_en : out STD_LOGIC;
           R57_en : out STD_LOGIC;
           R58_en : out STD_LOGIC;
           R59_en : out STD_LOGIC;
           R6_en : out STD_LOGIC;
           R60_en : out STD_LOGIC;
           R61_en : out STD_LOGIC;
           R62_en : out STD_LOGIC;
           R63_en : out STD_LOGIC;
           R64_en : out STD_LOGIC;
           R65_en : out STD_LOGIC;
           R66_en : out STD_LOGIC;
           R67_en : out STD_LOGIC;
           R68_en : out STD_LOGIC;
           R69_en : out STD_LOGIC;
           R7_en : out STD_LOGIC;
           R70_en : out STD_LOGIC;
           R71_en : out STD_LOGIC;
           R8_en : out STD_LOGIC;
           R9_en : out STD_LOGIC;
           A_en : out STD_LOGIC;
           A_wr : out STD_LOGIC;
           C_en : out STD_LOGIC;
           C_wr : out STD_LOGIC;
           W_en : out STD_LOGIC;
           W_wr : out STD_LOGIC;
           Mux_A_addr_sel : out STD_LOGIC_VECTOR(3 downto 0);
           Mux_Add_0_left_sel : out STD_LOGIC_VECTOR(3 downto 0);
           Mux_Add_0_right_sel : out STD_LOGIC_VECTOR(3 downto 0);
           Mux_C_addr_sel : out STD_LOGIC_VECTOR(3 downto 0);
           Mux_C_data_sel : out STD_LOGIC_VECTOR(3 downto 0);
           Mux_Mul_0_left_sel : out STD_LOGIC_VECTOR(3 downto 0);
           Mux_Mul_0_right_sel : out STD_LOGIC_VECTOR(3 downto 0);
           Mux_W_addr_sel : out STD_LOGIC_VECTOR(3 downto 0);
           state_out : out STD_LOGIC_VECTOR(4 downto 0));
end Controller;

architecture Behavioral of Controller is
    type state_type is (S0, S1, S2, S3, S4, S5, S6, S7, S8, S9, S10, S11, S12, S13, S14, S15, S_END);
    signal state : state_type := S0;
    function encode_state(s: state_type) return STD_LOGIC_VECTOR is
    begin
        case s is
            when S0 => return std_logic_vector(to_unsigned(0, 5));
            when S1 => return std_logic_vector(to_unsigned(1, 5));
            when S2 => return std_logic_vector(to_unsigned(2, 5));
            when S3 => return std_logic_vector(to_unsigned(3, 5));
            when S4 => return std_logic_vector(to_unsigned(4, 5));
            when S5 => return std_logic_vector(to_unsigned(5, 5));
            when S6 => return std_logic_vector(to_unsigned(6, 5));
            when S7 => return std_logic_vector(to_unsigned(7, 5));
            when S8 => return std_logic_vector(to_unsigned(8, 5));
            when S9 => return std_logic_vector(to_unsigned(9, 5));
            when S10 => return std_logic_vector(to_unsigned(10, 5));
            when S11 => return std_logic_vector(to_unsigned(11, 5));
            when S12 => return std_logic_vector(to_unsigned(12, 5));
            when S13 => return std_logic_vector(to_unsigned(13, 5));
            when S14 => return std_logic_vector(to_unsigned(14, 5));
            when S15 => return std_logic_vector(to_unsigned(15, 5));
            when S_END => return std_logic_vector(to_unsigned(16, 5));
        end case;
    end function;
begin

    process(clk, rst)
    begin
        if rst = '1' then state <= S0;
        elsif rising_edge(clk) then
            case state is
                when S0 => state <= S1;
                when S1 => state <= S2;
                when S2 => state <= S3;
                when S3 => state <= S4;
                when S4 => state <= S5;
                when S5 => state <= S6;
                when S6 => state <= S7;
                when S7 => state <= S8;
                when S8 => state <= S9;
                when S9 => state <= S10;
                when S10 => state <= S11;
                when S11 => state <= S12;
                when S12 => state <= S13;
                when S13 => state <= S14;
                when S14 => state <= S15;
                when S15 => state <= S_END;
                when others => state <= S_END;
            end case;
        end if;
    end process;

    state_out <= encode_state(state);

    process(state)
    begin
        R0_en <= '0';
        R1_en <= '0';
        R10_en <= '0';
        R11_en <= '0';
        R12_en <= '0';
        R13_en <= '0';
        R14_en <= '0';
        R15_en <= '0';
        R16_en <= '0';
        R17_en <= '0';
        R18_en <= '0';
        R19_en <= '0';
        R2_en <= '0';
        R20_en <= '0';
        R21_en <= '0';
        R22_en <= '0';
        R23_en <= '0';
        R24_en <= '0';
        R25_en <= '0';
        R26_en <= '0';
        R27_en <= '0';
        R28_en <= '0';
        R29_en <= '0';
        R3_en <= '0';
        R30_en <= '0';
        R31_en <= '0';
        R32_en <= '0';
        R33_en <= '0';
        R34_en <= '0';
        R35_en <= '0';
        R36_en <= '0';
        R37_en <= '0';
        R38_en <= '0';
        R39_en <= '0';
        R4_en <= '0';
        R40_en <= '0';
        R41_en <= '0';
        R42_en <= '0';
        R43_en <= '0';
        R44_en <= '0';
        R45_en <= '0';
        R46_en <= '0';
        R47_en <= '0';
        R48_en <= '0';
        R49_en <= '0';
        R5_en <= '0';
        R50_en <= '0';
        R51_en <= '0';
        R52_en <= '0';
        R53_en <= '0';
        R54_en <= '0';
        R55_en <= '0';
        R56_en <= '0';
        R57_en <= '0';
        R58_en <= '0';
        R59_en <= '0';
        R6_en <= '0';
        R60_en <= '0';
        R61_en <= '0';
        R62_en <= '0';
        R63_en <= '0';
        R64_en <= '0';
        R65_en <= '0';
        R66_en <= '0';
        R67_en <= '0';
        R68_en <= '0';
        R69_en <= '0';
        R7_en <= '0';
        R70_en <= '0';
        R71_en <= '0';
        R8_en <= '0';
        R9_en <= '0';
        A_en <= '0'; A_wr <= '0';
        C_en <= '0'; C_wr <= '0';
        W_en <= '0'; W_wr <= '0';
        Mux_A_addr_sel <= (others => '0');
        Mux_Add_0_left_sel <= (others => '0');
        Mux_Add_0_right_sel <= (others => '0');
        Mux_C_addr_sel <= (others => '0');
        Mux_C_data_sel <= (others => '0');
        Mux_Mul_0_left_sel <= (others => '0');
        Mux_Mul_0_right_sel <= (others => '0');
        Mux_W_addr_sel <= (others => '0');
        case state is
            when S0 =>
                R16_en <= '1';
                R0_en <= '1';
                R1_en <= '1';
                R4_en <= '1';
                R5_en <= '1';
                R10_en <= '1';
                R11_en <= '1';
                R34_en <= '1';
                R18_en <= '1';
                R19_en <= '1';
                R22_en <= '1';
                R23_en <= '1';
                R28_en <= '1';
                R29_en <= '1';
                R52_en <= '1';
                R36_en <= '1';
                R37_en <= '1';
                R40_en <= '1';
                R41_en <= '1';
                R46_en <= '1';
                R47_en <= '1';
                R70_en <= '1';
                R54_en <= '1';
                R55_en <= '1';
                R58_en <= '1';
                R59_en <= '1';
                R64_en <= '1';
                R65_en <= '1';
            when S1 =>
                R2_en <= '1';
                R3_en <= '1';
                A_en <= '1';
                W_en <= '1';
                Mux_A_addr_sel <= std_logic_vector(to_unsigned(0, 4));
                Mux_W_addr_sel <= std_logic_vector(to_unsigned(0, 4));
            when S2 =>
                R8_en <= '1';
                R6_en <= '1';
                R7_en <= '1';
                A_en <= '1';
                W_en <= '1';
                Mux_Mul_0_left_sel <= std_logic_vector(to_unsigned(0, 4));
                Mux_Mul_0_right_sel <= std_logic_vector(to_unsigned(0, 4));
                Mux_A_addr_sel <= std_logic_vector(to_unsigned(1, 4));
                Mux_W_addr_sel <= std_logic_vector(to_unsigned(1, 4));
            when S3 =>
                R9_en <= '1';
                R12_en <= '1';
                R13_en <= '1';
                A_en <= '1';
                W_en <= '1';
                Mux_Mul_0_left_sel <= std_logic_vector(to_unsigned(1, 4));
                Mux_Mul_0_right_sel <= std_logic_vector(to_unsigned(1, 4));
                Mux_A_addr_sel <= std_logic_vector(to_unsigned(2, 4));
                Mux_W_addr_sel <= std_logic_vector(to_unsigned(2, 4));
            when S4 =>
                R14_en <= '1';
                R15_en <= '1';
                R20_en <= '1';
                R21_en <= '1';
                A_en <= '1';
                W_en <= '1';
                Mux_Add_0_left_sel <= std_logic_vector(to_unsigned(0, 4));
                Mux_Add_0_right_sel <= std_logic_vector(to_unsigned(0, 4));
                Mux_Mul_0_left_sel <= std_logic_vector(to_unsigned(2, 4));
                Mux_Mul_0_right_sel <= std_logic_vector(to_unsigned(2, 4));
                Mux_A_addr_sel <= std_logic_vector(to_unsigned(3, 4));
                Mux_W_addr_sel <= std_logic_vector(to_unsigned(3, 4));
            when S5 =>
                R17_en <= '1';
                R26_en <= '1';
                R24_en <= '1';
                R25_en <= '1';
                A_en <= '1';
                W_en <= '1';
                Mux_Add_0_left_sel <= std_logic_vector(to_unsigned(1, 4));
                Mux_Add_0_right_sel <= std_logic_vector(to_unsigned(1, 4));
                Mux_Mul_0_left_sel <= std_logic_vector(to_unsigned(3, 4));
                Mux_Mul_0_right_sel <= std_logic_vector(to_unsigned(3, 4));
                Mux_A_addr_sel <= std_logic_vector(to_unsigned(4, 4));
                Mux_W_addr_sel <= std_logic_vector(to_unsigned(4, 4));
            when S6 =>
                R27_en <= '1';
                R30_en <= '1';
                R31_en <= '1';
                C_en <= '1';
                C_wr <= '1';
                A_en <= '1';
                W_en <= '1';
                Mux_C_addr_sel <= std_logic_vector(to_unsigned(0, 4));
                Mux_C_data_sel <= std_logic_vector(to_unsigned(0, 4));
                Mux_Mul_0_left_sel <= std_logic_vector(to_unsigned(4, 4));
                Mux_Mul_0_right_sel <= std_logic_vector(to_unsigned(4, 4));
                Mux_A_addr_sel <= std_logic_vector(to_unsigned(5, 4));
                Mux_W_addr_sel <= std_logic_vector(to_unsigned(5, 4));
            when S7 =>
                R32_en <= '1';
                R33_en <= '1';
                R38_en <= '1';
                R39_en <= '1';
                A_en <= '1';
                W_en <= '1';
                Mux_Add_0_left_sel <= std_logic_vector(to_unsigned(2, 4));
                Mux_Add_0_right_sel <= std_logic_vector(to_unsigned(2, 4));
                Mux_Mul_0_left_sel <= std_logic_vector(to_unsigned(5, 4));
                Mux_Mul_0_right_sel <= std_logic_vector(to_unsigned(5, 4));
                Mux_A_addr_sel <= std_logic_vector(to_unsigned(6, 4));
                Mux_W_addr_sel <= std_logic_vector(to_unsigned(6, 4));
            when S8 =>
                R35_en <= '1';
                R44_en <= '1';
                R42_en <= '1';
                R43_en <= '1';
                A_en <= '1';
                W_en <= '1';
                Mux_Add_0_left_sel <= std_logic_vector(to_unsigned(3, 4));
                Mux_Add_0_right_sel <= std_logic_vector(to_unsigned(3, 4));
                Mux_Mul_0_left_sel <= std_logic_vector(to_unsigned(6, 4));
                Mux_Mul_0_right_sel <= std_logic_vector(to_unsigned(6, 4));
                Mux_A_addr_sel <= std_logic_vector(to_unsigned(7, 4));
                Mux_W_addr_sel <= std_logic_vector(to_unsigned(7, 4));
            when S9 =>
                R45_en <= '1';
                R48_en <= '1';
                R49_en <= '1';
                C_en <= '1';
                C_wr <= '1';
                A_en <= '1';
                W_en <= '1';
                Mux_C_addr_sel <= std_logic_vector(to_unsigned(1, 4));
                Mux_C_data_sel <= std_logic_vector(to_unsigned(1, 4));
                Mux_Mul_0_left_sel <= std_logic_vector(to_unsigned(7, 4));
                Mux_Mul_0_right_sel <= std_logic_vector(to_unsigned(7, 4));
                Mux_A_addr_sel <= std_logic_vector(to_unsigned(8, 4));
                Mux_W_addr_sel <= std_logic_vector(to_unsigned(8, 4));
            when S10 =>
                R50_en <= '1';
                R51_en <= '1';
                R56_en <= '1';
                R57_en <= '1';
                A_en <= '1';
                W_en <= '1';
                Mux_Add_0_left_sel <= std_logic_vector(to_unsigned(4, 4));
                Mux_Add_0_right_sel <= std_logic_vector(to_unsigned(4, 4));
                Mux_Mul_0_left_sel <= std_logic_vector(to_unsigned(8, 4));
                Mux_Mul_0_right_sel <= std_logic_vector(to_unsigned(8, 4));
                Mux_A_addr_sel <= std_logic_vector(to_unsigned(9, 4));
                Mux_W_addr_sel <= std_logic_vector(to_unsigned(9, 4));
            when S11 =>
                R53_en <= '1';
                R62_en <= '1';
                R60_en <= '1';
                R61_en <= '1';
                A_en <= '1';
                W_en <= '1';
                Mux_Add_0_left_sel <= std_logic_vector(to_unsigned(5, 4));
                Mux_Add_0_right_sel <= std_logic_vector(to_unsigned(5, 4));
                Mux_Mul_0_left_sel <= std_logic_vector(to_unsigned(9, 4));
                Mux_Mul_0_right_sel <= std_logic_vector(to_unsigned(9, 4));
                Mux_A_addr_sel <= std_logic_vector(to_unsigned(10, 4));
                Mux_W_addr_sel <= std_logic_vector(to_unsigned(10, 4));
            when S12 =>
                R63_en <= '1';
                R66_en <= '1';
                R67_en <= '1';
                C_en <= '1';
                C_wr <= '1';
                A_en <= '1';
                W_en <= '1';
                Mux_C_addr_sel <= std_logic_vector(to_unsigned(2, 4));
                Mux_C_data_sel <= std_logic_vector(to_unsigned(2, 4));
                Mux_Mul_0_left_sel <= std_logic_vector(to_unsigned(10, 4));
                Mux_Mul_0_right_sel <= std_logic_vector(to_unsigned(10, 4));
                Mux_A_addr_sel <= std_logic_vector(to_unsigned(11, 4));
                Mux_W_addr_sel <= std_logic_vector(to_unsigned(11, 4));
            when S13 =>
                R68_en <= '1';
                R69_en <= '1';
                Mux_Add_0_left_sel <= std_logic_vector(to_unsigned(6, 4));
                Mux_Add_0_right_sel <= std_logic_vector(to_unsigned(6, 4));
                Mux_Mul_0_left_sel <= std_logic_vector(to_unsigned(11, 4));
                Mux_Mul_0_right_sel <= std_logic_vector(to_unsigned(11, 4));
            when S14 =>
                R71_en <= '1';
                Mux_Add_0_left_sel <= std_logic_vector(to_unsigned(7, 4));
                Mux_Add_0_right_sel <= std_logic_vector(to_unsigned(7, 4));
            when S15 =>
                C_en <= '1';
                C_wr <= '1';
                Mux_C_addr_sel <= std_logic_vector(to_unsigned(3, 4));
                Mux_C_data_sel <= std_logic_vector(to_unsigned(3, 4));
            when others => null;
        end case;
    end process;
end Behavioral;